library verilog;
use verilog.vl_types.all;
entity room_state is
end room_state;
