library verilog;
use verilog.vl_types.all;
entity lab04_02_sv_unit is
end lab04_02_sv_unit;
