library verilog;
use verilog.vl_types.all;
entity room_machine_sv_unit is
end room_machine_sv_unit;
