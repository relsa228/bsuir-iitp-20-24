package room_state;
typedef enum logic [3:0]{r_0, r_1, r_2, r_3, r_4, r_5, r_6, r_7} room_state_type;									
endpackage 